`timescale 1ns / 1ps 

module error1.v(clk, rst, );

input clk, rst;


endmodule
