`timescale 1ns / 1ps 

module m4(clk, rst, );

input clk, rst;


endmodule
