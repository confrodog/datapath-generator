`timescale 1ns / 1ps 

module error3.v(clk, rst, );

input clk, rst;


endmodule
