`timescale 1ns / 1ps 

module m5(clk, rst, );

input clk, rst;


endmodule
