`timescale 1ns / 1ps 

module error2.v(clk, rst, );

input clk, rst;


endmodule
